module uart_16550 ();

endmodule